`include "d_ff.v"

module tb_d_ff;

reg  d,clk, rst;
wire q;

d_ff dff (q, d, clk, rst); 
//Always at rising edge of clock display the signals
always @(posedge clk or negedge clk)begin
$display($time,"d=%b, clk=%b, rst=%b, q=%b\n", d, clk, rst, q);
end
//Module to generate clock with period 10 time units
initial 
begin
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
#5
clk=1;
#5
clk=0;
end

initial begin
d=0; rst=1;
#4
d=1; rst=0;
#50
d=1; rst=1;
#20
d=0; rst=0;
end
endmodule