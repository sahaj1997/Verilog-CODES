module ANDarray (Operation,Func,ALUOp1,ALUOp2);
input [3:0] Func;
input ALUOp1,ALUOp2;
output [2:0] Operation;


assign Op[0]= ;

assign Op[1]= ;

assign Op[3]= ;

endmodule